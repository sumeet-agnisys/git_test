
package hw_pkg;
    import uvm_pkg::*;
    import chip_name_regmem_pkg::*;
    import config_pkg::*;
    typedef enum {READ,WRITE} txn_kind;
        `include "uvm_macros.svh"

        //`include "agents/hardware_agent/hw_txn.svh"
        //`include "agents/hardware_agent/hw_adapter.svh"
        //`include "agents/hardware_agent/hw_driver.svh"
        //`include "agents/hardware_agent/hw_monitor.svh"
        //`include "agents/hardware_agent/hw_agent.svh"
    endpackage
