`define default_count         300 // Randomization repeated for 300 times.

`define reg_swRW_seq         `default_count // Randomization repeated 'default_count' for uvm_reg_swRW_seq
`define reg_swRO_seq         `default_count // Randomization repeated 'default_count' for uvm_reg_swRO_seq
`define reg_swWO_seq         `default_count // Randomization repeated 'default_count' for uvm_reg_swWO_seq
`define field_swRW_seq       `default_count // Randomization repeated 'default_count' for uvm_field_swRW_seq
`define field_swRO_seq       `default_count // Randomization repeated 'default_count' for uvm_field_swRO_seq
`define field_swWwtSE_seq    `default_count // Randomization repeated 'default_count' for uvm_field_swWwtSE_seq
`define field_swWO_seq       `default_count // Randomization repeated 'default_count' for uvm_field_swWO_seq
`define field_swRCRS_seq     `default_count // Randomization repeated 'default_count' for uvm_field_swRCRS_seq
`define field_swWRCWRS_seq   `default_count // Randomization repeated 'default_count' for uvm_field_swWRCWRS_seq
`define field_swWSRCWCRS_seq `default_count // Randomization repeated 'default_count' for uvm_field_swWSRCWCRS_seq
`define shadow_reg_seq       `default_count // Randomization repeated 'default_count' for shadow_reg_seq
`define alias_reg_seq       `default_count // Randomization repeated 'default_count' for alias_reg_seq
`define invalid_addr_seq       `default_count