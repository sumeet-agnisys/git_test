package seq_pkg;
 
    import arv_seq_pkg::*;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
    
	
	`include "seq_class.sv"
	
endpackage